`ifndef _my_params_h
`define _my_params_h
localparam OP_NOP = 4'd0;
localparam OP_MOV = 4'd1;
localparam OP_SWP = 4'd2;
localparam OP_SAV = 4'd3;
localparam OP_ADD = 4'd4;
localparam OP_SUB = 4'd5;
localparam OP_NEG = 4'd6;
localparam OP_JMP = 4'd7;
localparam OP_JEZ = 4'd8;
localparam OP_JNZ = 4'd9;
localparam OP_JGZ = 4'd10;
localparam OP_JLZ = 4'd11;
localparam OP_JRO = 4'd12;
`endif
