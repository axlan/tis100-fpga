`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/11/2020 05:34:23 PM
// Design Name: 
// Module Name: T21Node
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module t21_node(
        input clk,
        input reset,
        input signed [10:0] left_in_data,
        input signed left_in_ready,
        input signed [10:0] right_in_data,
        input signed right_in_ready,
        input signed [10:0] up_in_data,
        input signed up_in_ready,
        input signed [10:0] down_in_data,
        input signed down_in_ready,
        output signed [10:0] left_out_data,
        output signed left_out_ready,
        output signed [10:0] right_out_data,
        output signed right_out_ready,
        output signed [10:0] up_out_data,
        output signed up_out_ready,
        output signed [10:0] down_out_data,
        output signed down_out_ready
    );


    
    
    // alu alu_0()
    // instr_rom instr_rom_0()
    
    
    




endmodule
